localparam [31:0] BUILD_DATE = 32'h20200426;
localparam [31:0] BUILD_TIME = 32'h23163000;
