/*
Copyright (c) 2020 Chengdu JinZhiLi Technology Co., Ltd.
All rights reserved.
*/

parameter [7:0] VERSION_MAJOR = 8'd0;
parameter [7:0] VERSION_MINOR = 8'd9;
parameter [7:0] VERSION_PATCH = 8'd3;
parameter [7:0] VERSION_TWEAK = 8'd0;
