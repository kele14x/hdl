localparam [31:0] BUILD_DATE = 32'h20200423;
localparam [31:0] BUILD_TIME = 32'h10193300;
