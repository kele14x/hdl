/*
Copyright (c) 2019 Chengdu JinZhiLi Technology Co., Ltd.
All rights reserved.
*/

localparam [31:0] BUILD_DATE = 32'h20200630;
localparam [31:0] BUILD_TIME = 32'h09400000;
