localparam [31:0] BUILD_DATE = 32'h20200424;
localparam [31:0] BUILD_TIME = 32'h11173000;
