parameter [7:0] VERSION_MAJOR = 8'd0;
parameter [7:0] VERSION_MINOR = 8'd6;
parameter [7:0] VERSION_PATCH = 8'd0;
parameter [7:0] VERSION_TWEAK = 8'd1;
